//counter_tb.v

` timescale 1 ns / 1 ns

module tb_TOP_Counter();
  wire [7:0] CNT;
  reg [7:0] DATA;
  reg RST, CLK, LOAD, ENA;
  
  TOP_Counter UUT(CNT, DATA, CLK, RST, ENA, LOAD);
  //CLK Generator
  initial begin
    CLK = 1'b0;
    forever #10 CLK = ~CLK;
  end
  
  initial
    $monitorb("%d CLK = %b ENA = %b RST = %b CNT[7]= %b CNT[6]= %b CNT[5]= %b CNT[4]= %b CNT[3]= %b CNT[2]= %b CNT[1]= %b CNT[0]= %b",$time, CLK, ENA, RST, CNT[7], CNT[6], CNT[5], CNT[4], CNT[3], CNT[2],CNT[1], CNT[0]);

  initial begin
    $vcdpluson;
    // Demonstrates Asynchronous Reset
    #10 $display ("\n Demonstrates Asynchronous Reset\n"); RST =
    1'b0;
    // Counter initiates
    #20 $display ("\n Counter initiates\n"); ENA = 1'b1; RST = 1'b1;
    LOAD = 1'b0;
    // After 8 there is parallel load of 250
    #200 $display ("\n After 8 there is parallel load of 250\n"); ENA
    = 1'b1; LOAD = 1'b1; DATA = 8'd250;
    //Starts counting from 250 and rolls over
    #20 $display ("\n Starts counting from 250\n"); LOAD = 1'b0;
    //Reset overrides Load
    #140 $display ("\n Reset overrides load\n"); LOAD = 1'b1; RST =
    1'b0;
    // Reset overrides increment
    #40 $display ("\n Reset overrides increment\n"); LOAD = 1'b0; ENA
    = 1'b1; RST = 1'b0; DATA = 8'd10;
    #60 ENA = 1'b1; RST = 1'b1; LOAD = 1'b0;
    //Enable low for Load
    #140 $display ("\n Enable low for Load\n"); LOAD = 1'b1; ENA =
    1'b0;
    // Enable low for increment
    #40 $display ("\n Enable low for increment \n"); LOAD = 1'b0; ENA
    = 1'b0; DATA = 8'd200;
    //#40 $stop;
    #40 $finish;
  end
endmodule